package pyst;
  import uvm_pkg::*;

  `include "param.sv"
  `include "argument.sv"
  `include "packet.sv"
  `include "service_subscriber.sv"
  `include "service.sv"
endpackage : pyst
