package rp_component;
  import uvm_pkg::*;
  `include "common.sv"
endpackage